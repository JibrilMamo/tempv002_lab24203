parameter LW = 6'b100011 ; 
parameter SW = 6'b101011 ;
parameter no_op = 32'b0000000_0000000_0000000_0000000 ;
parameter ALUop = 6'b0 ;
parameter CINDC = 54 ;
parameter BEQINIT = 55 ;
//C:\Users\Kartik\Documents\solution_lab2_fall_2023\solution
string filename="/export/scratch/users/ramkr004/solution_lab2_fall_2023/solution/testing_path/regs.dat";
string filename1="/export/scratch/users/ramkr004/solution_lab2_fall_2023/solution/testing_path/dmem.dat";
string filename2="/export/scratch/users/ramkr004/solution_lab2_fall_2023/solution/testing_path/imem.dat";
string filename3="/export/scratch/users/ramkr004/solution_lab2_fall_2023/solution/testing_path/mem_result.dat";
string filename4="/export/scratch/users/ramkr004/solution_lab2_fall_2023/solution/testing_path/regs_result.dat";